CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 0 5 200 9
1968 106 3792 997
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
1968 106 3792 997
177209362 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 587 204 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 457 159 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 540 138 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 535 98 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 SR Flip-Flop~
219 773 134 0 4 9
0 2 16 3 17
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
2 U5
25 -34 39 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
9 Inverter~
13 700 101 0 2 22
0 2 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7734 0 0
0
0
9 2-In AND~
219 677 253 0 3 22
0 9 10 2
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
9 2-In NOR~
219 758 237 0 3 22
0 7 8 10
0
0 0 624 180
6 74LS02
-21 -24 21 -16
3 U4A
7 -25 28 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3747 0 0
0
0
9 2-In AND~
219 767 276 0 3 22
0 5 6 9
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3549 0 0
0
0
14 Logic Display~
6 734 158 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
12 Hex Display~
7 848 132 0 18 19
10 5 7 6 8 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9325 0 0
0
0
7 74LS169
9 660 176 0 14 29
0 14 15 13 2 2 12 2 4 3
11 8 6 7 5
0
0 0 13040 0
6 74F169
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
22
1 0 2 0 0 8192 0 5 0 0 5 4
784 81
784 76
699 76
699 75
9 3 3 0 0 12416 0 12 5 0 0 5
692 149
722 149
722 142
766 142
766 135
4 0 2 0 0 0 0 12 0 0 5 4
628 185
616 185
616 181
604 181
8 2 4 0 0 8320 0 12 6 0 0 3
698 140
703 140
703 119
1 3 2 0 0 12416 0 6 7 0 0 5
703 83
703 75
604 75
604 253
650 253
0 1 5 0 0 4096 0 0 9 22 0 3
834 212
834 285
785 285
0 2 6 0 0 4096 0 0 9 20 0 3
823 194
823 267
785 267
0 1 7 0 0 4096 0 0 8 21 0 3
809 203
809 246
783 246
0 2 8 0 0 4096 0 0 8 19 0 3
800 185
800 228
783 228
3 1 9 0 0 4224 0 9 7 0 0 4
740 276
708 276
708 262
695 262
3 2 10 0 0 4224 0 8 7 0 0 4
731 237
708 237
708 244
695 244
1 10 11 0 0 4224 0 10 12 0 0 2
734 176
698 176
7 0 2 0 0 0 0 12 0 0 5 2
628 212
604 212
5 0 2 0 0 0 0 12 0 0 5 4
628 194
612 194
612 186
604 186
1 6 12 0 0 8320 0 1 12 0 0 3
599 204
599 203
628 203
3 1 13 0 0 4224 0 12 2 0 0 4
628 158
483 158
483 159
469 159
1 1 14 0 0 4224 0 12 4 0 0 4
622 140
558 140
558 98
547 98
2 1 15 0 0 4224 0 12 3 0 0 4
622 149
561 149
561 138
552 138
4 11 8 0 0 8320 0 11 12 0 0 3
839 156
839 185
692 185
3 12 6 0 0 8320 0 11 12 0 0 3
845 156
845 194
692 194
13 2 7 0 0 4224 0 12 11 0 0 3
692 203
851 203
851 156
1 14 5 0 0 8320 0 11 12 0 0 3
857 156
857 212
692 212
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
