CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
177209362 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 134 290 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 199 110 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
9 Inverter~
13 300 598 0 2 22
0 10 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3618 0 0
0
0
9 Inverter~
13 305 515 0 2 22
0 8 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
6153 0 0
0
0
14 Logic Display~
6 858 552 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
8 4-In OR~
219 732 569 0 5 22
0 6 5 3 4 2
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 -1969888268
65 0 0 0 2 1 5 0
1 U
7734 0 0
0
0
9 2-In AND~
219 508 655 0 3 22
0 8 7 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9914 0 0
0
0
9 2-In AND~
219 508 608 0 3 22
0 9 7 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3747 0 0
0
0
9 2-In AND~
219 510 559 0 3 22
0 9 7 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
9 2-In AND~
219 512 499 0 3 22
0 9 10 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7931 0 0
0
0
8 3-In OR~
219 673 302 0 4 22
0 14 13 12 11
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 3 0
1 U
9325 0 0
0
0
14 Logic Display~
6 835 295 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
9 2-In AND~
219 513 418 0 3 22
0 8 15 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3834 0 0
0
0
9 2-In AND~
219 521 308 0 3 22
0 16 15 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3363 0 0
0
0
9 2-In AND~
219 512 193 0 3 22
0 16 10 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7668 0 0
0
0
9 Inverter~
13 319 327 0 2 22
0 10 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4718 0 0
0
0
9 Inverter~
13 397 185 0 2 22
0 8 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3874 0 0
0
0
27
5 1 2 0 0 8320 0 6 5 0 0 3
765 569
765 570
858 570
3 3 3 0 0 4224 0 6 8 0 0 4
715 574
588 574
588 608
529 608
4 3 4 0 0 12416 0 6 7 0 0 4
715 583
663 583
663 655
529 655
2 3 5 0 0 4224 0 6 9 0 0 4
715 565
543 565
543 559
531 559
3 1 6 0 0 4224 0 10 6 0 0 4
533 499
646 499
646 556
715 556
2 0 7 0 0 4096 0 8 0 0 7 2
484 617
357 617
0 2 7 0 0 0 0 0 7 10 0 3
357 598
357 664
484 664
0 1 8 0 0 8192 0 0 7 15 0 3
238 515
238 646
484 646
0 1 9 0 0 4096 0 0 8 11 0 3
461 548
461 599
484 599
2 2 7 0 0 12416 0 3 9 0 0 4
321 598
357 598
357 568
486 568
0 1 9 0 0 4096 0 0 9 14 0 3
461 490
461 550
486 550
0 2 10 0 0 4096 0 0 10 13 0 4
266 537
423 537
423 508
488 508
0 1 10 0 0 4224 0 0 3 23 0 3
266 327
266 598
285 598
2 1 9 0 0 4224 0 4 10 0 0 4
326 515
411 515
411 490
488 490
0 1 8 0 0 4224 0 0 4 27 0 3
238 185
238 515
290 515
4 1 11 0 0 4224 0 11 12 0 0 4
706 302
803 302
803 313
835 313
3 3 12 0 0 4224 0 13 11 0 0 4
534 418
650 418
650 311
660 311
3 2 13 0 0 4224 0 14 11 0 0 4
542 308
635 308
635 302
661 302
3 1 14 0 0 4224 0 15 11 0 0 4
533 193
642 193
642 293
660 293
1 2 10 0 0 128 0 16 15 0 0 3
304 327
304 202
488 202
2 2 15 0 0 8192 0 16 13 0 0 3
340 327
340 427
489 427
2 2 15 0 0 8320 0 16 14 0 0 3
340 327
340 317
497 317
1 1 10 0 0 0 0 1 16 0 0 4
146 290
263 290
263 327
304 327
2 1 16 0 0 4224 0 17 14 0 0 3
418 185
418 299
497 299
1 1 8 0 0 128 0 17 13 0 0 3
382 185
382 409
489 409
2 1 16 0 0 0 0 17 15 0 0 3
418 185
418 184
488 184
1 1 8 0 0 0 0 2 17 0 0 4
211 110
238 110
238 185
382 185
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
