CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 816 1872 1004
193986578 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 92 61 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
5 SCOPE
12 622 187 0 1 11
0 2
0
0 0 57584 0
4 TP11
-14 -4 14 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4441 0 0
0
0
9 2-In AND~
219 750 304 0 3 22
0 4 3 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3618 0 0
0
0
10 2-In NAND~
219 885 313 0 3 22
0 6 5 2
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6153 0 0
0
0
12 Hex Display~
7 553 28 0 16 19
10 3 4 5 7 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5394 0 0
0
0
5 SCOPE
12 1158 132 0 1 11
0 7
0
0 0 57584 0
4 TP10
-14 -4 14 4
2 U7
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 831 130 0 1 11
0 5
0
0 0 57584 0
3 TP9
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 469 129 0 1 11
0 4
0
0 0 57584 0
3 TP7
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 189 139 0 1 11
0 3
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 86 148 0 1 11
0 9
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
14 Logic Display~
6 1187 125 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
6 JK RN~
219 1111 159 0 6 22
0 8 5 8 2 10 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
8903 0 0
0
0
6 JK RN~
219 782 158 0 6 22
0 8 4 8 2 11 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3834 0 0
0
0
14 Logic Display~
6 858 124 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
6 JK RN~
219 427 157 0 6 22
0 8 3 8 2 12 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
7668 0 0
0
0
14 Logic Display~
6 503 123 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
6 JK RN~
219 146 167 0 6 22
0 8 9 8 2 13 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
3874 0 0
0
0
14 Logic Display~
6 222 133 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
7 Pulser~
4 55 170 0 10 12
0 14 15 9 16 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3789 0 0
0
0
34
1 0 2 0 0 4096 0 2 0 0 21 2
622 199
622 198
2 0 3 0 0 4224 0 3 0 0 31 3
726 313
199 313
199 151
1 0 4 0 0 4224 0 3 0 0 30 3
726 295
458 295
458 141
0 2 5 0 0 4096 0 0 4 29 0 3
818 142
818 322
861 322
3 1 6 0 0 4224 0 3 4 0 0 2
771 304
861 304
3 0 2 0 0 8192 0 4 0 0 20 3
912 313
919 313
919 198
2 1 5 0 0 4096 0 12 14 0 0 3
1080 151
858 151
858 142
2 0 4 0 0 128 0 13 0 0 30 3
751 150
497 150
497 141
1 2 3 0 0 0 0 18 15 0 0 3
222 151
222 149
396 149
4 0 7 0 0 8320 0 5 0 0 28 4
544 52
544 108
1175 108
1175 143
3 0 5 0 0 8320 0 5 0 0 29 4
550 52
550 88
848 88
848 142
1 0 3 0 0 128 0 5 0 0 31 4
562 52
562 98
207 98
207 151
2 0 4 0 0 128 0 5 0 0 30 4
556 52
556 78
489 78
489 141
1 0 4 0 0 0 0 8 0 0 30 2
469 141
469 141
0 0 8 0 0 4096 0 0 0 27 33 4
367 58
132 58
132 103
92 103
1 0 7 0 0 0 0 6 0 0 28 2
1158 144
1158 143
1 0 5 0 0 0 0 7 0 0 29 2
831 142
831 142
1 0 3 0 0 0 0 9 0 0 31 2
189 151
189 151
1 0 9 0 0 4096 0 10 0 0 34 2
86 160
86 159
0 4 2 0 0 4096 0 0 12 21 0 3
781 198
1111 198
1111 190
0 4 2 0 0 4224 0 0 13 22 0 3
426 198
782 198
782 189
4 4 2 0 0 0 0 17 15 0 0 3
146 198
427 198
427 188
1 0 8 0 0 0 0 12 0 0 25 2
1087 142
1046 142
1 0 8 0 0 0 0 13 0 0 25 2
758 141
721 141
3 3 8 0 0 12416 0 13 12 0 0 6
758 159
721 159
721 58
1046 58
1046 160
1087 160
1 0 8 0 0 0 0 15 0 0 27 2
403 140
366 140
0 3 8 0 0 4224 0 0 15 25 0 4
721 58
366 58
366 158
403 158
6 1 7 0 0 128 0 12 11 0 0 3
1135 142
1135 143
1187 143
6 1 5 0 0 128 0 13 14 0 0 3
806 141
806 142
858 142
6 1 4 0 0 128 0 15 16 0 0 3
451 140
451 141
503 141
6 1 3 0 0 128 0 17 18 0 0 3
170 150
170 151
222 151
1 0 8 0 0 0 0 17 0 0 33 2
122 150
92 150
1 3 8 0 0 128 0 1 17 0 0 3
92 73
92 168
122 168
3 2 9 0 0 8320 0 19 17 0 0 3
79 161
79 159
115 159
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
