CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
440 210 4 200 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
0 71 1920 1040
177209362 256
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 693 468 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 603 378 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 720 360 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
9 Inverter~
13 828 504 0 2 22
0 5 9
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
6153 0 0
0
0
9 Inverter~
13 819 504 0 2 22
0 6 10
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
5394 0 0
0
0
12 SPDT Switch~
164 639 414 0 3 11
0 13 12 13
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7734 0 0
0
0
13 SR Flip-Flop~
219 1089 432 0 4 9
0 11 4 16 21
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
9 Inverter~
13 891 603 0 2 22
0 17 11
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3747 0 0
0
0
9 Inverter~
13 828 603 0 2 22
0 2 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3549 0 0
0
0
9 Inverter~
13 891 504 0 2 22
0 5 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
7931 0 0
0
0
9 Inverter~
13 864 504 0 2 22
0 8 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9325 0 0
0
0
10 4-In NAND~
219 886 549 0 5 22
0 7 18 6 19 17
0
0 0 624 270
6 74LS20
-21 -28 21 -20
3 U3B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
8903 0 0
0
0
10 4-In NAND~
219 828 549 0 5 22
0 7 9 10 8 2
0
0 0 624 270
6 74LS20
-21 -28 21 -20
3 U3A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 -151122343
65 0 0 0 2 1 2 0
1 U
3834 0 0
0
0
9 2-In NOR~
219 990 405 0 3 22
0 4 11 15
0
0 0 624 180
6 74LS02
-21 -24 21 -16
3 U2A
7 -25 28 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3363 0 0
0
0
7 Pulser~
4 576 432 0 10 12
0 22 23 13 24 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7668 0 0
0
0
12 Hex Display~
7 918 315 0 18 19
10 7 5 6 8 0 0 0 0 0
0 1 0 0 1 1 1 0 12
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4718 0 0
0
0
7 74LS169
9 774 441 0 14 29
0 20 20 13 2 2 3 2 15 16
25 8 6 5 7
0
0 0 13040 0
6 74F169
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
33
7 0 2 0 0 4096 0 17 0 0 3 2
742 477
731 477
5 0 2 0 0 0 0 17 0 0 3 2
742 459
731 459
0 4 2 0 0 8320 0 0 17 21 0 4
829 581
731 581
731 450
742 450
1 6 3 0 0 4224 0 1 17 0 0 2
705 468
742 468
0 1 4 0 0 4096 0 0 14 12 0 2
1055 414
1015 414
1 0 5 0 0 4096 0 4 0 0 31 2
831 486
831 468
1 0 6 0 0 4096 0 5 0 0 32 2
822 486
822 459
1 0 7 0 0 4096 0 13 0 0 30 2
842 524
842 477
4 0 8 0 0 4096 0 13 0 0 33 2
815 524
815 450
2 2 9 0 0 4224 0 4 13 0 0 3
831 522
831 524
833 524
2 3 10 0 0 4224 0 5 13 0 0 3
822 522
822 524
824 524
2 2 4 0 0 12416 0 9 7 0 0 5
831 621
831 639
1055 639
1055 414
1065 414
0 2 11 0 0 4224 0 0 8 14 0 3
1035 396
1035 621
894 621
1 2 11 0 0 0 0 7 14 0 0 2
1065 396
1015 396
1 2 12 0 0 8320 0 2 6 0 0 6
615 378
620 378
620 405
617 405
617 410
622 410
1 3 13 0 0 4224 0 6 17 0 0 4
656 414
728 414
728 423
742 423
3 3 13 0 0 4224 14 15 6 0 0 4
600 423
614 423
614 418
622 418
3 8 15 0 0 4224 0 14 17 0 0 2
963 405
812 405
3 9 16 0 0 12416 0 7 17 0 0 6
1119 414
1156 414
1156 353
826 353
826 414
806 414
5 1 17 0 0 4224 0 12 8 0 0 3
887 575
887 585
894 585
5 1 2 0 0 128 0 13 9 0 0 3
829 575
829 585
831 585
0 1 7 0 0 0 0 0 12 30 0 3
906 477
906 524
900 524
0 1 5 0 0 0 0 0 10 31 0 2
894 468
894 486
0 3 6 0 0 4096 0 0 12 32 0 3
879 459
879 524
882 524
0 1 8 0 0 0 0 0 11 33 0 2
867 450
867 486
2 2 18 0 0 8320 0 10 12 0 0 3
894 522
894 524
891 524
2 4 19 0 0 8320 0 11 12 0 0 3
867 522
867 524
873 524
1 1 20 0 0 8320 0 17 3 0 0 6
736 405
732 405
732 370
738 370
738 360
732 360
2 1 20 0 0 0 0 17 17 0 0 2
736 414
736 405
1 14 7 0 0 4224 0 16 17 0 0 3
927 339
927 477
806 477
2 13 5 0 0 4224 0 16 17 0 0 3
921 339
921 468
806 468
3 12 6 0 0 4224 0 16 17 0 0 3
915 339
915 459
806 459
11 4 8 0 0 8320 0 17 16 0 0 3
806 450
909 450
909 339
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
