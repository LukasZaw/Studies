CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 9 200 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
0 71 1920 1040
177209362 256
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 414 162 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 225 162 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
9 2-In AND~
219 333 279 0 3 22
0 4 3 2
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3618 0 0
0
0
9 3-In AND~
219 522 252 0 4 22
0 5 6 7 4
0
0 0 624 270
6 74LS11
-21 -28 21 -20
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
6153 0 0
0
0
14 Logic Display~
6 279 90 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
7 Pulser~
4 378 288 0 10 12
0 15 16 8 17 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7734 0 0
0
0
12 Hex Display~
7 540 81 0 18 19
10 5 6 7 10 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9914 0 0
0
0
6 74LS90
107 459 189 0 10 21
0 9 9 2 2 8 5 10 7 6
5
0
0 0 13040 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
12 Hex Display~
7 333 90 0 16 19
10 11 12 13 3 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3549 0 0
0
0
6 74LS90
107 270 189 0 10 21
0 14 14 2 2 10 11 3 13 12
11
0
0 0 13040 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
26
3 4 2 0 0 12416 0 3 8 0 0 5
331 302
331 331
416 331
416 189
427 189
3 0 2 0 0 0 0 3 0 0 24 4
331 302
217 302
217 184
238 184
0 2 3 0 0 4224 0 0 3 22 0 2
322 162
322 257
4 1 4 0 0 8320 0 4 3 0 0 6
520 275
520 279
412 279
412 252
340 252
340 257
0 1 5 0 0 4096 0 0 4 14 0 2
529 216
529 230
0 2 6 0 0 4096 0 0 4 15 0 2
520 198
520 230
0 3 7 0 0 4096 0 0 4 16 0 3
503 180
503 230
511 230
5 3 8 0 0 8320 0 8 6 0 0 3
421 207
402 207
402 279
1 0 3 0 0 0 0 5 0 0 22 4
279 108
279 134
309 134
309 162
3 4 2 0 0 128 0 8 8 0 0 2
427 180
427 189
2 1 9 0 0 8320 0 8 1 0 0 3
427 171
426 171
426 162
1 1 9 0 0 0 0 1 8 0 0 2
426 162
427 162
0 5 10 0 0 8320 0 0 10 17 0 5
497 162
497 250
221 250
221 207
232 207
1 10 5 0 0 4224 0 7 8 0 0 3
549 105
549 216
491 216
2 9 6 0 0 4224 0 7 8 0 0 3
543 105
543 198
491 198
3 8 7 0 0 4224 0 7 8 0 0 3
537 105
537 180
491 180
7 4 10 0 0 0 0 8 7 0 0 3
491 162
531 162
531 105
6 10 5 0 0 0 0 8 8 0 0 4
421 216
421 227
491 227
491 216
1 10 11 0 0 4224 0 9 10 0 0 3
342 114
342 216
302 216
2 9 12 0 0 4224 0 9 10 0 0 3
336 114
336 198
302 198
3 8 13 0 0 4224 0 9 10 0 0 3
330 114
330 180
302 180
7 4 3 0 0 128 0 10 9 0 0 3
302 162
324 162
324 114
2 1 14 0 0 4224 0 10 10 0 0 2
238 171
238 162
4 3 2 0 0 128 0 10 10 0 0 2
238 189
238 180
1 1 14 0 0 0 0 2 10 0 0 2
237 162
238 162
6 10 11 0 0 128 0 10 10 0 0 4
232 216
232 232
302 232
302 216
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
