CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 0 10 200 9
1968 106 3792 997
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
1968 106 3792 997
177209362 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 571 319 0 1 11
0 2
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
12 Hex Display~
7 763 62 0 16 19
10 3 4 12 13 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
4441 0 0
0
0
12 Hex Display~
7 627 56 0 16 19
10 8 7 6 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3618 0 0
0
0
14 Logic Display~
6 694 311 0 1 2
10 9
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
9 4-In AND~
219 638 151 0 5 22
0 5 6 7 8 10
0
0 0 624 270
6 74LS21
-21 -28 21 -20
3 U4A
19 -4 40 4
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 -417962061
65 0 0 0 2 1 2 0
1 U
5394 0 0
0
0
9 2-In AND~
219 673 238 0 3 22
0 11 10 9
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7734 0 0
0
0
9 2-In AND~
219 705 197 0 3 22
0 3 4 11
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9914 0 0
0
0
6 74LS93
109 762 187 0 8 17
0 9 9 5 3 14 15 4 3
0
0 0 13040 90
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
6 74LS93
109 565 188 0 8 17
0 9 9 2 8 5 6 7 8
0
0 0 13040 90
6 74LS93
-21 -35 21 -27
2 U1
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
25
0 1 2 0 0 8192 0 0 1 20 0 3
570 279
572 279
572 306
8 1 3 0 0 4096 0 8 2 0 0 4
776 153
776 94
772 94
772 86
7 2 4 0 0 4096 0 8 2 0 0 4
767 153
767 94
766 94
766 86
0 4 5 0 0 4096 0 0 3 25 0 5
552 136
614 136
614 88
618 88
618 80
0 3 6 0 0 4096 0 0 3 13 0 5
561 127
614 127
614 88
624 88
624 80
0 2 7 0 0 4096 0 0 3 14 0 5
570 127
614 127
614 88
630 88
630 80
0 1 8 0 0 8192 0 0 3 15 0 5
579 136
614 136
614 88
636 88
636 80
0 1 9 0 0 4096 0 0 4 16 0 2
694 265
694 297
1 8 3 0 0 8192 0 7 8 0 0 4
712 175
712 145
776 145
776 153
2 7 4 0 0 12416 0 7 8 0 0 5
694 175
693 175
693 145
767 145
767 153
5 0 10 0 0 4224 0 5 0 0 19 2
636 174
636 223
0 1 5 0 0 4096 0 0 5 25 0 3
552 121
649 121
649 129
6 2 6 0 0 8320 0 9 5 0 0 4
561 154
561 121
640 121
640 129
7 3 7 0 0 8320 0 9 5 0 0 4
570 154
570 121
631 121
631 129
8 4 8 0 0 0 0 9 5 0 0 5
579 154
579 121
623 121
623 129
622 129
0 0 9 0 0 8192 0 0 0 17 21 4
664 261
664 265
754 265
754 217
0 3 9 0 0 8320 0 0 6 22 0 3
557 218
557 261
671 261
3 1 11 0 0 8320 0 7 6 0 0 3
703 220
703 216
680 216
2 0 10 0 0 0 0 6 0 0 0 3
662 216
662 223
635 223
3 0 2 0 0 4224 0 9 0 0 0 3
570 224
570 279
549 279
1 2 9 0 0 0 0 8 8 0 0 2
749 217
758 217
1 2 9 0 0 0 0 9 9 0 0 2
552 218
561 218
8 4 8 0 0 12416 0 9 9 0 0 6
579 154
579 150
594 150
594 232
579 232
579 224
8 4 3 0 0 12416 0 8 8 0 0 6
776 153
776 149
822 149
822 250
776 250
776 223
5 3 5 0 0 8320 0 9 8 0 0 6
552 154
552 101
800 101
800 235
767 235
767 223
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
