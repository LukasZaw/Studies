CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 171 538 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 467 345 0 1 11
0 26
0
0 0 21360 90
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 238 346 0 1 11
0 25
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 431 339 0 1 11
0 27
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 201 347 0 1 11
0 28
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 904 311 0 1 11
0 32
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 1134 303 0 1 11
0 31
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 70 436 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
14 Logic Display~
6 1189 137 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 1175 137 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 1160 137 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 1142 141 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 966 136 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 946 137 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 926 135 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 908 138 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
13 SR Flip-Flop~
219 266 548 0 4 9
0 20 19 21 33
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
12 Hex Display~
7 456 120 0 18 19
10 12 14 15 11 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6671 0 0
0
0
12 Hex Display~
7 238 128 0 18 19
10 13 16 17 18 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3789 0 0
0
0
9 2-In AND~
219 237 438 0 3 22
0 22 21 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4871 0 0
0
0
12 SPDT Switch~
164 157 433 0 3 11
0 22 24 22
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3750 0 0
0
0
6 74LS90
107 466 277 0 10 21
0 27 27 26 26 10 12 11 15 14
12
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U5
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
6 74LS90
107 238 286 0 10 21
0 28 28 25 25 11 13 18 17 16
13
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U4
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
6 74LS90
107 941 250 0 10 21
0 32 32 30 30 10 3 9 4 8
3
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U2
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
6 74LS90
107 1169 241 0 10 21
0 31 31 29 29 10 2 5 7 6
2
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U1
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
9 2-In AND~
219 1050 230 0 3 22
0 4 3 30
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5950 0 0
0
0
9 2-In AND~
219 1299 231 0 3 22
0 5 2 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5670 0 0
0
0
9 2-In AND~
219 1252 391 0 3 22
0 30 29 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6828 0 0
0
0
14 Logic Display~
6 1273 373 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
7 Pulser~
4 67 504 0 10 12
0 34 35 22 36 0 0 5 5 5
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8365 0 0
0
0
53
0 6 2 0 0 4096 0 0 25 6 0 4
1232 199
1232 281
1196 281
1196 273
0 6 3 0 0 4224 0 0 24 4 0 4
1004 199
1004 290
968 290
968 282
0 1 4 0 0 4224 0 0 26 13 0 3
926 193
1057 193
1057 208
0 2 3 0 0 0 0 0 26 11 0 3
966 199
1039 199
1039 208
0 1 5 0 0 4224 0 0 27 10 0 3
1142 192
1306 192
1306 209
0 2 2 0 0 8320 0 0 27 7 0 4
1195 195
1195 199
1288 199
1288 209
1 10 2 0 0 0 0 9 25 0 0 4
1189 155
1189 195
1196 195
1196 203
9 1 6 0 0 4224 0 25 10 0 0 4
1178 203
1178 163
1175 163
1175 155
1 8 7 0 0 4224 0 11 25 0 0 2
1160 155
1160 203
7 1 5 0 0 0 0 25 12 0 0 2
1142 203
1142 159
1 10 3 0 0 0 0 13 24 0 0 4
966 154
966 204
968 204
968 212
9 1 8 0 0 4224 0 24 14 0 0 4
950 212
950 163
946 163
946 155
1 8 4 0 0 0 0 15 24 0 0 4
926 153
926 204
932 204
932 212
7 1 9 0 0 4224 0 24 16 0 0 4
914 212
914 164
908 164
908 156
0 0 10 0 0 8320 0 0 0 31 16 4
959 384
959 433
483 433
483 438
3 5 10 0 0 0 0 20 22 0 0 3
258 438
484 438
484 309
0 5 11 0 0 4224 0 0 23 23 0 5
439 230
280 230
280 326
256 326
256 318
0 6 12 0 0 12288 0 0 22 20 0 6
493 231
493 235
508 235
508 317
493 317
493 309
0 6 13 0 0 12288 0 0 23 24 0 6
265 240
265 244
280 244
280 326
265 326
265 318
1 10 12 0 0 4224 0 18 22 0 0 4
465 144
465 231
493 231
493 239
9 2 14 0 0 4224 0 22 18 0 0 4
475 239
475 152
459 152
459 144
3 8 15 0 0 4224 0 18 22 0 0 4
453 144
453 231
457 231
457 239
7 4 11 0 0 0 0 22 18 0 0 4
439 239
439 152
447 152
447 144
1 10 13 0 0 4224 0 19 23 0 0 4
247 152
247 240
265 240
265 248
9 2 16 0 0 4224 0 23 19 0 0 4
247 248
247 160
241 160
241 152
3 8 17 0 0 4224 0 19 23 0 0 4
235 152
235 240
229 240
229 248
7 4 18 0 0 4224 0 23 19 0 0 4
211 248
211 160
229 160
229 152
1 2 19 0 0 4224 0 1 17 0 0 4
183 538
234 538
234 530
242 530
3 1 20 0 0 12416 0 28 17 0 0 6
1273 391
1285 391
1285 498
234 498
234 512
242 512
3 2 21 0 0 12416 0 17 20 0 0 6
296 530
300 530
300 458
205 458
205 447
213 447
5 5 10 0 0 0 0 25 24 0 0 4
1187 273
1187 384
959 384
959 282
1 1 22 0 0 4224 0 21 20 0 0 4
174 433
205 433
205 429
213 429
3 3 22 0 0 8320 23 21 30 0 0 4
140 437
105 437
105 495
91 495
2 1 24 0 0 4224 0 21 8 0 0 4
140 429
91 429
91 436
82 436
1 4 25 0 0 12416 0 3 23 0 0 4
239 333
239 326
238 326
238 312
1 3 26 0 0 4224 0 2 22 0 0 4
468 332
468 317
457 317
457 303
4 3 25 0 0 16 0 23 23 0 0 2
238 312
229 312
3 4 26 0 0 16 0 22 22 0 0 2
457 303
466 303
1 2 27 0 0 8336 0 4 22 0 0 4
432 326
432 317
448 317
448 303
1 1 27 0 0 16 0 4 22 0 0 4
432 326
432 317
439 317
439 303
2 1 28 0 0 8336 0 23 5 0 0 4
220 312
220 327
202 327
202 334
1 1 28 0 0 16 0 23 5 0 0 4
211 312
211 327
202 327
202 334
1 3 20 0 0 0 0 29 28 0 0 2
1273 391
1273 391
0 2 29 0 0 4096 0 0 28 47 0 3
1220 277
1220 400
1228 400
0 1 30 0 0 8320 0 0 28 46 0 4
1035 290
1035 344
1228 344
1228 382
3 4 30 0 0 0 0 26 24 0 0 4
1048 253
1048 290
941 290
941 276
4 3 29 0 0 8320 0 25 27 0 0 4
1169 267
1169 277
1297 277
1297 254
4 3 30 0 0 0 0 24 24 0 0 2
941 276
932 276
3 4 29 0 0 0 0 25 25 0 0 2
1160 267
1169 267
1 2 31 0 0 8320 0 7 25 0 0 4
1135 290
1135 281
1151 281
1151 267
1 1 31 0 0 0 0 7 25 0 0 4
1135 290
1135 281
1142 281
1142 267
2 1 32 0 0 8320 0 24 6 0 0 4
923 276
923 291
905 291
905 298
1 1 32 0 0 0 0 24 6 0 0 4
914 276
914 291
905 291
905 298
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
