CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 190 1 200 9
-1920 150 0 1119
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
-1920 873 0 1119
193986578 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 559 379 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 493 356 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 497 307 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 487 252 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 491 135 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5394 0 0
0
0
5 SCOPE
12 716 562 0 1 11
0 2
0
0 0 57584 0
3 TP4
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 550 538 0 1 11
0 3
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 375 529 0 1 11
0 4
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
14 Logic Display~
6 731 524 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
12 D Flip-Flop~
219 657 577 0 4 9
0 6 2 6 5
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 578 559 0 3 22
0 3 5 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 402 550 0 3 22
0 4 7 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8903 0 0
0
0
12 D Flip-Flop~
219 481 568 0 4 9
0 8 3 8 7
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
14 Logic Display~
6 548 415 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
12 D Flip-Flop~
219 486 476 0 4 9
0 10 4 10 9
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
14 Logic Display~
6 620 301 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
6 JK RN~
219 560 338 0 6 22
0 13 4 12 14 21 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3874 0 0
0
0
14 Logic Display~
6 695 149 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
9 2-In AND~
219 559 238 0 3 22
0 20 18 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3789 0 0
0
0
9 2-In AND~
219 570 160 0 3 22
0 19 20 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4871 0 0
0
0
13 SR Flip-Flop~
219 628 210 0 4 9
0 17 16 22 15
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
7 Pulser~
4 323 188 0 10 12
0 23 24 20 4 0 0 5 5 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8778 0 0
0
0
27
1 0 2 0 0 0 0 6 0 0 4 2
716 574
716 574
1 0 3 0 0 0 0 7 0 0 5 2
550 550
550 550
1 0 4 0 0 0 0 8 0 0 9 2
375 541
375 541
0 1 2 0 0 8320 0 0 9 8 0 4
623 559
623 574
731 574
731 542
0 1 3 0 0 8320 0 0 11 12 0 5
447 550
447 564
536 564
536 550
562 550
4 2 5 0 0 8320 0 10 11 0 0 5
681 541
681 585
554 585
554 568
562 568
1 3 6 0 0 8320 0 10 10 0 0 5
633 541
633 522
693 522
693 559
687 559
2 3 2 0 0 0 0 10 11 0 0 2
633 559
611 559
1 0 4 0 0 8192 0 12 0 0 13 3
386 541
358 541
358 458
4 2 7 0 0 8320 0 13 12 0 0 5
505 532
505 576
378 576
378 559
386 559
1 3 8 0 0 8320 0 13 13 0 0 5
457 532
457 513
517 513
517 550
511 550
2 3 3 0 0 0 0 13 12 0 0 2
457 550
435 550
2 0 4 0 0 8192 0 15 0 0 17 4
462 458
358 458
358 329
353 329
4 1 9 0 0 4224 0 15 14 0 0 3
510 440
548 440
548 433
1 3 10 0 0 12416 0 15 15 0 0 6
462 440
458 440
458 473
524 473
524 458
516 458
6 1 11 0 0 4224 0 17 16 0 0 5
584 321
608 321
608 327
620 327
620 319
4 2 4 0 0 8320 0 22 17 0 0 3
353 188
353 330
529 330
1 3 12 0 0 8320 0 2 17 0 0 4
505 356
521 356
521 339
536 339
1 1 13 0 0 12416 0 3 17 0 0 4
509 307
521 307
521 321
536 321
1 4 14 0 0 4224 0 1 17 0 0 2
560 366
560 369
4 1 15 0 0 4224 0 21 18 0 0 3
652 174
695 174
695 167
3 2 16 0 0 8320 0 19 21 0 0 4
580 238
596 238
596 192
604 192
3 1 17 0 0 8320 0 20 21 0 0 4
591 160
596 160
596 174
604 174
1 2 18 0 0 4224 0 4 19 0 0 4
499 252
524 252
524 247
535 247
1 1 19 0 0 4224 0 5 20 0 0 4
503 135
526 135
526 151
546 151
3 0 20 0 0 4224 0 22 0 0 27 2
347 179
524 179
2 1 20 0 0 128 0 20 19 0 0 4
546 169
524 169
524 229
535 229
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
