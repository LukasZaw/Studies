CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 113 288 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 184 87 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
12 Hex Display~
7 717 29 0 18 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3618 0 0
0
0
6 JK RN~
219 1269 232 0 6 22
0 9 7 9 6 11 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 6 0
1 U
6153 0 0
0
0
6 JK RN~
219 907 223 0 6 22
0 10 7 10 6 12 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 5 0
1 U
5394 0 0
0
0
6 JK RN~
219 547 219 0 6 22
0 5 7 5 6 13 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 5 0
1 U
7734 0 0
0
0
6 JK RN~
219 259 215 0 6 22
0 8 7 8 6 14 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 4 0
1 U
9914 0 0
0
0
5 SCOPE
12 1358 203 0 1 11
0 2
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 993 196 0 1 11
0 3
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 634 156 0 1 11
0 4
0
0 0 57584 270
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 371 186 0 1 11
0 5
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9325 0 0
0
0
14 Logic Display~
6 963 190 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 601 184 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 325 181 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 1467 127 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
7 Pulser~
4 85 202 0 10 12
0 15 16 7 17 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4718 0 0
0
0
9 2-In AND~
219 1092 102 0 3 22
0 10 3 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3874 0 0
0
0
9 2-In AND~
219 784 107 0 3 22
0 4 5 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
41
4 0 2 0 0 8320 0 3 0 0 37 4
708 53
708 73
1388 73
1388 215
3 0 3 0 0 8320 0 3 0 0 21 4
714 53
714 60
1026 60
1026 207
2 0 4 0 0 4096 0 3 0 0 28 2
720 53
720 98
1 0 5 0 0 8320 0 3 0 0 29 4
726 53
726 88
410 88
410 198
4 0 6 0 0 4096 0 4 0 0 13 2
1269 263
1269 265
2 0 7 0 0 0 0 4 0 0 38 2
1238 224
1238 224
4 0 6 0 0 0 0 5 0 0 24 2
907 254
907 254
2 0 7 0 0 4096 0 5 0 0 39 2
876 215
876 216
4 0 6 0 0 0 0 6 0 0 23 2
547 250
548 250
2 0 7 0 0 0 0 6 0 0 40 2
516 211
516 211
4 0 6 0 0 0 0 7 0 0 22 2
259 246
258 246
2 0 7 0 0 0 0 7 0 0 41 2
228 207
228 207
0 0 6 0 0 8192 0 0 0 25 0 3
1269 265
1267 265
1267 257
1 0 2 0 0 0 0 8 0 0 37 2
1358 215
1358 215
1 0 3 0 0 0 0 9 0 0 21 2
993 208
993 207
1 0 4 0 0 0 0 10 0 0 28 2
625 159
626 159
1 0 5 0 0 0 0 11 0 0 29 2
371 198
371 198
1 0 3 0 0 0 0 12 0 0 21 2
963 208
963 207
1 0 4 0 0 0 0 13 0 0 28 2
601 202
601 202
1 0 5 0 0 0 0 14 0 0 29 2
325 199
325 198
6 2 3 0 0 0 0 5 17 0 0 5
931 206
931 207
1060 207
1060 111
1068 111
0 0 6 0 0 4096 0 0 0 0 25 2
258 240
258 288
0 0 6 0 0 0 0 0 0 0 25 2
548 244
548 288
0 0 6 0 0 0 0 0 0 0 25 2
907 249
907 288
1 0 6 0 0 4224 0 1 0 0 0 4
125 288
1269 288
1269 257
1267 257
0 2 5 0 0 0 0 0 18 29 0 3
496 202
496 116
760 116
3 0 5 0 0 0 0 6 0 0 29 3
523 220
506 220
506 202
6 1 4 0 0 12416 0 6 18 0 0 4
571 202
626 202
626 98
760 98
6 1 5 0 0 0 0 7 6 0 0 4
283 198
458 198
458 202
523 202
0 3 8 0 0 8192 0 0 7 31 0 3
184 196
184 216
235 216
1 1 8 0 0 4224 0 2 7 0 0 3
184 99
184 198
235 198
1 0 9 0 0 4096 0 4 0 0 33 2
1245 215
1228 215
3 3 9 0 0 8320 0 17 4 0 0 4
1113 102
1228 102
1228 233
1245 233
0 3 10 0 0 4096 0 0 5 35 0 4
865 207
865 225
883 225
883 224
0 1 10 0 0 4096 0 0 5 36 0 4
847 107
847 207
883 207
883 206
3 1 10 0 0 4224 0 18 17 0 0 4
805 107
1043 107
1043 93
1068 93
6 1 2 0 0 0 0 4 15 0 0 3
1293 215
1467 215
1467 145
0 0 7 0 0 4224 0 0 0 39 0 4
848 266
1214 266
1214 224
1243 224
0 0 7 0 0 0 0 0 0 40 0 4
483 266
848 266
848 216
883 216
0 0 7 0 0 0 0 0 0 41 0 5
154 207
154 266
484 266
484 211
524 211
3 0 7 0 0 0 0 16 0 0 0 4
109 193
154 193
154 207
234 207
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
