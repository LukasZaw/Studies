CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 816 1872 1004
193986578 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 166 407 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 600 211 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 92 61 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
9 Inverter~
13 804 350 0 2 22
0 2 14
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
6153 0 0
0
0
9 Inverter~
13 473 342 0 2 22
0 2 17
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
5394 0 0
0
0
9 Inverter~
13 175 338 0 2 22
0 2 20
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
7734 0 0
0
0
8 2-In OR~
219 906 346 0 3 22
0 12 13 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9914 0 0
0
0
8 2-In OR~
219 572 336 0 3 22
0 16 15 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3747 0 0
0
0
8 2-In OR~
219 287 329 0 3 22
0 19 18 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3549 0 0
0
0
9 2-In AND~
219 847 399 0 3 22
0 5 2 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7931 0 0
0
0
9 2-In AND~
219 841 305 0 3 22
0 4 14 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9325 0 0
0
0
9 2-In AND~
219 519 385 0 3 22
0 8 2 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8903 0 0
0
0
9 2-In AND~
219 518 300 0 3 22
0 7 17 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3834 0 0
0
0
9 2-In AND~
219 223 369 0 3 22
0 11 2 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3363 0 0
0
0
9 2-In AND~
219 220 299 0 3 22
0 10 20 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7668 0 0
0
0
12 Hex Display~
7 553 28 0 18 19
10 10 7 4 21 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4718 0 0
0
0
5 SCOPE
12 1158 132 0 1 11
0 21
0
0 0 57584 0
4 TP10
-14 -4 14 4
2 U7
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3874 0 0
0
0
5 SCOPE
12 831 130 0 1 11
0 4
0
0 0 57584 0
3 TP9
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6671 0 0
0
0
5 SCOPE
12 469 129 0 1 11
0 7
0
0 0 57584 0
3 TP7
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3789 0 0
0
0
5 SCOPE
12 189 139 0 1 11
0 10
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4871 0 0
0
0
5 SCOPE
12 86 148 0 1 11
0 23
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3750 0 0
0
0
14 Logic Display~
6 1187 125 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
6 JK RN~
219 1111 159 0 6 22
0 22 3 22 24 25 21
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
538 0 0
0
0
6 JK RN~
219 782 158 0 6 22
0 22 6 22 24 5 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
6843 0 0
0
0
14 Logic Display~
6 858 124 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
6 JK RN~
219 427 157 0 6 22
0 22 9 22 24 8 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
5950 0 0
0
0
14 Logic Display~
6 503 123 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5670 0 0
0
0
6 JK RN~
219 146 167 0 6 22
0 22 23 22 24 11 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
6828 0 0
0
0
14 Logic Display~
6 222 133 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
7 Pulser~
4 55 170 0 10 12
0 26 27 23 28 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8365 0 0
0
0
50
1 0 2 0 0 4096 0 1 0 0 2 2
178 407
178 408
0 0 2 0 0 4096 0 0 0 3 24 3
477 408
178 408
178 378
0 0 2 0 0 4224 0 0 0 15 20 3
808 408
476 408
476 394
3 2 3 0 0 4224 0 7 23 0 0 3
939 346
939 151
1080 151
1 0 4 0 0 4096 0 11 0 0 45 2
817 296
817 142
5 1 5 0 0 12416 0 24 10 0 0 5
812 159
812 236
753 236
753 390
823 390
3 2 6 0 0 8320 0 8 24 0 0 4
605 336
666 336
666 150
751 150
1 0 7 0 0 8336 0 13 0 0 46 3
494 291
464 291
464 141
1 5 8 0 0 8320 0 12 26 0 0 3
495 376
457 376
457 158
3 2 9 0 0 4224 0 9 26 0 0 3
320 329
320 149
396 149
0 1 10 0 0 4096 0 0 15 47 0 3
178 151
178 290
196 290
5 1 11 0 0 16512 0 28 14 0 0 6
176 168
188 168
188 254
134 254
134 360
199 360
3 1 12 0 0 4224 0 11 7 0 0 3
862 305
862 337
893 337
3 2 13 0 0 4224 0 10 7 0 0 3
868 399
868 355
893 355
2 1 2 0 0 128 0 10 4 0 0 3
823 408
807 408
807 368
2 2 14 0 0 4224 0 4 11 0 0 3
807 332
807 314
817 314
2 3 15 0 0 8320 0 8 12 0 0 4
559 345
546 345
546 385
540 385
3 1 16 0 0 4224 0 13 8 0 0 3
539 300
539 327
559 327
2 2 17 0 0 8320 0 5 13 0 0 3
476 324
476 309
494 309
2 1 2 0 0 128 0 12 5 0 0 3
495 394
476 394
476 360
3 2 18 0 0 4224 0 14 9 0 0 3
244 369
244 338
274 338
3 1 19 0 0 8320 0 15 9 0 0 4
241 299
258 299
258 320
274 320
2 2 20 0 0 8320 0 6 15 0 0 3
178 320
178 308
196 308
2 1 2 0 0 128 0 14 6 0 0 3
199 378
178 378
178 356
4 0 21 0 0 8320 0 16 0 0 44 4
544 52
544 108
1175 108
1175 143
3 0 4 0 0 8320 0 16 0 0 45 4
550 52
550 88
848 88
848 142
1 0 10 0 0 8320 0 16 0 0 47 4
562 52
562 98
207 98
207 151
2 0 7 0 0 128 0 16 0 0 46 4
556 52
556 78
489 78
489 141
1 0 7 0 0 0 0 19 0 0 46 2
469 141
469 141
0 0 22 0 0 4096 0 0 0 43 49 4
367 58
132 58
132 103
92 103
1 0 21 0 0 0 0 17 0 0 44 2
1158 144
1158 143
1 0 4 0 0 0 0 18 0 0 45 2
831 142
831 142
1 0 10 0 0 0 0 20 0 0 47 2
189 151
189 151
1 0 23 0 0 4096 0 21 0 0 50 2
86 160
86 159
1 0 24 0 0 0 0 2 0 0 37 2
601 198
601 198
0 4 24 0 0 4096 0 0 23 37 0 3
781 198
1111 198
1111 190
0 4 24 0 0 4224 0 0 24 38 0 3
426 198
782 198
782 189
4 4 24 0 0 0 0 28 26 0 0 3
146 198
427 198
427 188
1 0 22 0 0 0 0 23 0 0 41 2
1087 142
1046 142
1 0 22 0 0 0 0 24 0 0 41 2
758 141
721 141
3 3 22 0 0 12416 0 24 23 0 0 6
758 159
721 159
721 58
1046 58
1046 160
1087 160
1 0 22 0 0 0 0 26 0 0 43 2
403 140
366 140
0 3 22 0 0 4224 0 0 26 41 0 4
721 58
366 58
366 158
403 158
6 1 21 0 0 128 0 23 22 0 0 3
1135 142
1135 143
1187 143
6 1 4 0 0 128 0 24 25 0 0 3
806 141
806 142
858 142
6 1 7 0 0 128 0 26 27 0 0 3
451 140
451 141
503 141
6 1 10 0 0 128 0 28 29 0 0 3
170 150
170 151
222 151
1 0 22 0 0 0 0 28 0 0 49 2
122 150
92 150
1 3 22 0 0 128 0 3 28 0 0 3
92 73
92 168
122 168
3 2 23 0 0 8320 0 30 28 0 0 3
79 161
79 159
115 159
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
