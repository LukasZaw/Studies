CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 120 9 200 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
0 71 1920 1040
177209362 256
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 405 315 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 603 315 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
10 2-In NAND~
219 747 405 0 3 22
0 3 4 2
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U4A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3618 0 0
0
0
9 2-In AND~
219 783 324 0 3 22
0 7 8 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6153 0 0
0
0
9 2-In AND~
219 549 324 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5394 0 0
0
0
9 2-In AND~
219 585 387 0 3 22
0 10 2 9
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U3A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7734 0 0
0
0
7 Pulser~
4 522 423 0 10 12
0 17 18 10 19 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9914 0 0
0
0
12 Hex Display~
7 513 216 0 18 19
10 14 5 6 16 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3747 0 0
0
0
12 Hex Display~
7 747 225 0 18 19
10 8 7 15 13 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3549 0 0
0
0
6 74LS93
109 648 324 0 8 17
0 12 12 9 8 13 15 7 8
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
6 74LS93
109 450 324 0 8 17
0 11 11 13 14 16 6 5 14
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
24
3 2 2 0 0 8320 0 3 6 0 0 4
748 431
748 435
593 435
593 408
3 1 3 0 0 12416 0 4 3 0 0 5
804 324
808 324
808 372
757 372
757 380
3 2 4 0 0 12416 0 5 3 0 0 5
570 324
603 324
603 372
739 372
739 380
2 0 5 0 0 8192 0 5 0 0 22 3
525 333
525 330
516 330
1 0 6 0 0 4096 0 5 0 0 23 2
525 315
510 315
1 0 7 0 0 8192 0 4 0 0 18 3
759 315
759 312
750 312
2 0 8 0 0 4096 0 4 0 0 17 3
759 333
759 338
756 338
3 3 9 0 0 4224 0 6 10 0 0 3
584 363
584 333
610 333
1 3 10 0 0 8320 0 6 7 0 0 3
575 408
575 414
546 414
1 2 11 0 0 4224 0 11 11 0 0 2
418 315
418 324
1 2 12 0 0 4224 0 10 10 0 0 2
616 315
616 324
1 1 11 0 0 0 0 1 11 0 0 2
417 315
418 315
1 1 12 0 0 0 0 2 10 0 0 2
615 315
616 315
0 3 13 0 0 8320 0 0 11 20 0 5
687 315
687 259
382 259
382 333
412 333
4 0 14 0 0 12288 0 11 0 0 21 5
412 342
408 342
408 357
491 357
491 342
4 0 8 0 0 12288 0 10 0 0 17 5
610 342
606 342
606 357
686 357
686 342
1 8 8 0 0 4224 0 9 10 0 0 3
756 249
756 342
680 342
2 7 7 0 0 4224 0 9 10 0 0 3
750 249
750 333
680 333
3 6 15 0 0 4224 0 9 10 0 0 3
744 249
744 324
680 324
4 5 13 0 0 0 0 9 10 0 0 3
738 249
738 315
680 315
1 8 14 0 0 4224 0 8 11 0 0 3
522 240
522 342
482 342
2 7 5 0 0 4224 0 8 11 0 0 3
516 240
516 333
482 333
3 6 6 0 0 4224 0 8 11 0 0 3
510 240
510 324
482 324
4 5 16 0 0 4224 0 8 11 0 0 3
504 240
504 315
482 315
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
