CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
811 114 2635 1012
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
811 849 2635 1012
193986578 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 173 152 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 927 248 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 85 407 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
5 SCOPE
12 987 143 0 1 11
0 2
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 751 144 0 1 11
0 3
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 554 157 0 1 11
0 4
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 330 153 0 1 11
0 5
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 116 318 0 1 11
0 6
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
14 Logic Display~
6 940 136 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 715 138 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 501 153 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 285 148 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
9 Inverter~
13 125 182 0 2 22
0 7 11
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3834 0 0
0
0
6 JK RN~
219 867 173 0 6 22
0 3 6 8 12 13 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3363 0 0
0
0
6 JK RN~
219 664 186 0 6 22
0 4 6 9 12 8 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
7668 0 0
0
0
6 JK RN~
219 452 183 0 6 22
0 5 6 10 12 9 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
4718 0 0
0
0
6 JK RN~
219 234 182 0 6 22
0 7 6 11 12 10 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3874 0 0
0
0
7 Pulser~
4 67 330 0 10 12
0 14 15 16 6 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6671 0 0
0
0
28
1 0 2 0 0 4096 0 4 0 0 6 2
987 155
987 154
1 0 3 0 0 0 0 5 0 0 12 2
751 156
751 156
1 0 4 0 0 0 0 6 0 0 15 2
554 169
554 169
1 0 5 0 0 0 0 7 0 0 16 2
330 165
330 165
1 0 6 0 0 4096 0 8 0 0 21 2
116 330
116 329
1 0 2 0 0 4224 0 9 0 0 0 2
940 154
993 154
6 1 2 0 0 0 0 14 9 0 0 3
891 156
891 154
940 154
1 0 3 0 0 0 0 10 0 0 12 2
715 156
715 156
1 0 4 0 0 4096 0 11 0 0 15 2
501 171
501 169
1 0 5 0 0 4096 0 12 0 0 16 2
285 166
285 165
1 0 7 0 0 0 0 1 0 0 19 2
173 164
173 164
1 6 3 0 0 4224 0 14 15 0 0 3
843 156
688 156
688 169
5 3 8 0 0 4224 0 15 14 0 0 3
694 187
843 187
843 174
3 5 9 0 0 4224 0 15 16 0 0 3
640 187
482 187
482 184
6 1 4 0 0 8320 0 16 15 0 0 3
476 166
476 169
640 169
1 6 5 0 0 8320 0 16 17 0 0 3
428 166
428 165
258 165
5 3 10 0 0 8320 0 17 16 0 0 3
264 183
264 184
428 184
2 3 11 0 0 4224 0 13 17 0 0 4
128 200
203 200
203 183
210 183
1 1 7 0 0 8320 0 17 13 0 0 3
210 165
210 164
128 164
1 0 6 0 0 8192 0 3 0 0 21 3
97 407
136 407
136 329
4 0 6 0 0 8192 0 18 0 0 28 3
97 330
97 329
179 329
1 0 12 0 0 8192 0 2 0 0 25 3
913 248
913 228
866 228
4 0 12 0 0 0 0 15 0 0 25 2
664 217
664 228
4 0 12 0 0 0 0 16 0 0 25 2
452 214
452 228
4 4 12 0 0 8320 0 17 14 0 0 4
234 213
234 228
867 228
867 204
2 0 6 0 0 8192 0 15 0 0 28 3
633 178
628 178
628 329
2 0 6 0 0 8192 0 16 0 0 28 3
421 175
414 175
414 329
2 2 6 0 0 12416 0 14 17 0 0 6
836 165
825 165
825 329
179 329
179 174
203 174
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
