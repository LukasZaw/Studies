CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
814 114 2638 1012
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
814 114 2638 1012
177209362 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 70 451 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 185 598 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 326 198 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 127 271 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
5 SCOPE
12 480 34 0 1 11
0 3
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 411 34 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 355 34 0 1 11
0 2
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
14 Logic Display~
6 1046 384 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 647 385 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 324 386 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
9 2-In AND~
219 140 388 0 3 22
0 8 9 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9325 0 0
0
0
9 Inverter~
13 380 170 0 2 22
0 13 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
8903 0 0
0
0
8 2-In OR~
219 836 405 0 3 22
0 16 15 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3834 0 0
0
0
9 3-In AND~
219 746 446 0 4 22
0 17 12 13 15
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 5 0
1 U
3363 0 0
0
0
9 3-In AND~
219 746 370 0 4 22
0 11 2 4 16
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
7668 0 0
0
0
8 2-In OR~
219 495 412 0 3 22
0 20 19 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4718 0 0
0
0
9 2-In AND~
219 424 457 0 3 22
0 12 13 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3874 0 0
0
0
9 2-In AND~
219 423 369 0 3 22
0 11 2 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
7 Pulser~
4 53 389 0 10 12
0 21 22 8 23 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3789 0 0
0
0
12 Hex Display~
7 183 28 0 18 19
10 2 4 3 5 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4871 0 0
0
0
14 Logic Display~
6 1687 323 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3750 0 0
0
0
6 JK RN~
219 1395 421 0 6 22
0 25 26 27 28 29 30
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
8778 0 0
0
0
6 JK RN~
219 1000 419 0 6 22
0 14 7 14 10 31 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
538 0 0
0
0
6 JK RN~
219 608 419 0 6 22
0 18 7 18 10 17 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
6843 0 0
0
0
6 JK RN~
219 288 419 0 6 22
0 6 7 6 10 12 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3136 0 0
0
0
43
0 1 2 0 0 4224 0 0 0 42 12 2
320 402
320 66
1 3 3 0 0 4096 0 5 0 0 12 2
480 46
480 66
1 2 4 0 0 4096 0 6 0 0 12 2
411 46
411 66
1 1 2 0 0 0 0 7 0 0 12 2
355 46
355 66
1 3 3 0 0 8320 0 8 0 0 12 5
1046 402
1066 402
1066 99
940 99
940 66
6 1 3 0 0 0 0 23 8 0 0 2
1024 402
1046 402
0 2 4 0 0 4224 0 0 0 37 12 2
637 402
637 66
4 4 5 0 0 4224 0 20 0 0 12 2
174 52
174 66
3 3 3 0 0 0 0 20 0 0 12 2
180 52
180 66
2 2 4 0 0 0 0 20 0 0 12 2
186 52
186 66
1 1 2 0 0 0 0 20 0 0 12 2
192 52
192 66
-6369869 0 1 0 0 4256 0 0 0 0 0 2
75 66
976 66
1 0 4 0 0 0 0 9 0 0 37 2
647 403
647 402
1 0 2 0 0 0 0 10 0 0 42 2
324 404
324 402
0 1 6 0 0 4224 0 0 4 16 0 3
247 402
247 271
139 271
3 1 6 0 0 0 0 25 25 0 0 4
264 420
247 420
247 402
264 402
3 0 7 0 0 8192 0 11 0 0 21 4
161 388
189 388
189 442
241 442
3 1 8 0 0 8320 0 19 11 0 0 3
77 380
77 379
116 379
2 1 9 0 0 8320 0 11 1 0 0 4
116 397
99 397
99 451
82 451
0 2 7 0 0 4224 0 0 23 21 0 4
567 573
958 573
958 411
969 411
2 2 7 0 0 0 0 25 24 0 0 6
257 411
241 411
241 573
568 573
568 411
577 411
4 0 10 0 0 8192 0 23 0 0 24 3
1000 450
1000 598
604 598
4 0 10 0 0 0 0 25 0 0 24 2
288 450
288 598
1 4 10 0 0 4224 0 2 24 0 0 3
197 598
608 598
608 450
0 2 2 0 0 0 0 0 15 42 0 5
374 378
374 304
692 304
692 370
722 370
1 2 11 0 0 8192 0 18 12 0 0 3
399 360
401 360
401 170
2 1 11 0 0 4224 0 12 15 0 0 4
401 170
717 170
717 361
722 361
0 2 12 0 0 8320 0 0 14 43 0 5
367 420
367 489
685 489
685 446
722 446
2 0 13 0 0 4096 0 17 0 0 30 2
400 466
344 466
0 3 13 0 0 4224 0 0 14 31 0 5
344 197
344 558
705 558
705 455
722 455
1 1 13 0 0 0 0 12 3 0 0 4
365 170
344 170
344 198
338 198
3 0 14 0 0 4224 0 13 0 0 33 2
869 405
949 405
3 1 14 0 0 0 0 23 23 0 0 4
976 420
949 420
949 402
976 402
2 4 15 0 0 4224 0 13 14 0 0 4
823 414
786 414
786 446
767 446
4 1 16 0 0 12416 0 15 13 0 0 4
767 370
787 370
787 396
823 396
1 5 17 0 0 4224 0 14 24 0 0 4
722 437
675 437
675 420
638 420
6 3 4 0 0 0 0 24 15 0 0 4
632 402
676 402
676 379
722 379
0 3 18 0 0 8320 0 0 24 39 0 3
556 412
556 420
584 420
3 1 18 0 0 0 0 16 24 0 0 4
528 412
556 412
556 402
584 402
2 3 19 0 0 8320 0 16 17 0 0 4
482 421
454 421
454 457
445 457
3 1 20 0 0 8320 0 18 16 0 0 4
444 369
454 369
454 403
482 403
6 2 2 0 0 0 0 25 18 0 0 4
312 402
374 402
374 378
399 378
1 5 12 0 0 0 0 17 25 0 0 4
400 448
373 448
373 420
318 420
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
